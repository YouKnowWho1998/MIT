module pipe(
    input wire sys_clk 
    input 
)